/* lu.v
 * LU module implementation, calculate logic
 * with different input modes
 */
`include "def.v"


